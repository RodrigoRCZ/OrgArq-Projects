module decoder1035(input c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11,output s);

    assign s = c1 & ~c2 & ~c3 & ~c4 & ~c5 & ~c6 & ~c7 & c8 & ~c9 & c10 & c11;

endmodule